library verilog;
use verilog.vl_types.all;
entity ParamCounter_tb is
end ParamCounter_tb;
