library verilog;
use verilog.vl_types.all;
entity Factorial_tb is
end Factorial_tb;
