library verilog;
use verilog.vl_types.all;
entity AlwaysTest_tb is
end AlwaysTest_tb;
