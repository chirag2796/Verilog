library verilog;
use verilog.vl_types.all;
entity DFlipFlopWithEnable_tb is
end DFlipFlopWithEnable_tb;
