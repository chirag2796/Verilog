library verilog;
use verilog.vl_types.all;
entity DFlipFlopWithReset_tb is
end DFlipFlopWithReset_tb;
