library verilog;
use verilog.vl_types.all;
entity ClkGen1 is
    port(
        clk             : out    vl_logic
    );
end ClkGen1;
