library verilog;
use verilog.vl_types.all;
entity HalfAdderOp_tb is
end HalfAdderOp_tb;
