library verilog;
use verilog.vl_types.all;
entity \NOT\ is
    port(
        a               : in     vl_logic;
        o               : out    vl_logic
    );
end \NOT\;
