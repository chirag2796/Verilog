library verilog;
use verilog.vl_types.all;
entity MUX_4TO1 is
    port(
        i0              : in     vl_logic;
        i1              : in     vl_logic;
        i2              : in     vl_logic;
        i3              : in     vl_logic;
        s0              : in     vl_logic;
        s1              : in     vl_logic;
        o               : out    vl_logic
    );
end MUX_4TO1;
