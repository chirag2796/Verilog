library verilog;
use verilog.vl_types.all;
entity ClkForever is
    port(
        clk             : out    vl_logic
    );
end ClkForever;
