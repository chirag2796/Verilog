library verilog;
use verilog.vl_types.all;
entity reduction_op_tb is
end reduction_op_tb;
