library verilog;
use verilog.vl_types.all;
entity for_example is
end for_example;
