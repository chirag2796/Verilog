library verilog;
use verilog.vl_types.all;
entity Multiply is
    port(
        a               : in     vl_logic_vector(7 downto 0);
        b               : in     vl_logic_vector(7 downto 0);
        ans             : out    vl_logic_vector(15 downto 0)
    );
end Multiply;
