library verilog;
use verilog.vl_types.all;
entity Bh_HalfAdder_tb is
end Bh_HalfAdder_tb;
