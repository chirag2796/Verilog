library verilog;
use verilog.vl_types.all;
entity halfsubtractor_tb is
end halfsubtractor_tb;
