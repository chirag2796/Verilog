library verilog;
use verilog.vl_types.all;
entity bit_counter_tb is
end bit_counter_tb;
