library verilog;
use verilog.vl_types.all;
entity mux_4to1_tb is
end mux_4to1_tb;
