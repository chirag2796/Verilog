library verilog;
use verilog.vl_types.all;
entity DLatchWithoutResetEnable_tb is
end DLatchWithoutResetEnable_tb;
