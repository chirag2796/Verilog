library verilog;
use verilog.vl_types.all;
entity while_example_tb is
end while_example_tb;
