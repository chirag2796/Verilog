library verilog;
use verilog.vl_types.all;
entity RepeatMemory is
end RepeatMemory;
