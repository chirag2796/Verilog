library verilog;
use verilog.vl_types.all;
entity DLatchWithResetEnable_tb is
end DLatchWithResetEnable_tb;
