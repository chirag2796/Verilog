library verilog;
use verilog.vl_types.all;
entity DLatchWithReset_tb is
end DLatchWithReset_tb;
