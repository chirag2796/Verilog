library verilog;
use verilog.vl_types.all;
entity DLatchWithEnable_tb is
end DLatchWithEnable_tb;
