library verilog;
use verilog.vl_types.all;
entity arithmetic_op_tb is
end arithmetic_op_tb;
