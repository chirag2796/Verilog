library verilog;
use verilog.vl_types.all;
entity Decoder2to4Op_tb is
end Decoder2to4Op_tb;
