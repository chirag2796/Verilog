library verilog;
use verilog.vl_types.all;
entity FunctionCalling_tb is
end FunctionCalling_tb;
