library verilog;
use verilog.vl_types.all;
entity RepeatCounter is
end RepeatCounter;
