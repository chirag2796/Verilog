library verilog;
use verilog.vl_types.all;
entity DFlipFlopWithResetEnable_tb is
end DFlipFlopWithResetEnable_tb;
