library verilog;
use verilog.vl_types.all;
entity DFlipFlopWithoutResetEnable_tb is
end DFlipFlopWithoutResetEnable_tb;
