library verilog;
use verilog.vl_types.all;
entity not_tb is
end not_tb;
