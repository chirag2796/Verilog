library verilog;
use verilog.vl_types.all;
entity Multiply_tb is
end Multiply_tb;
