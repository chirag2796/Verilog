library verilog;
use verilog.vl_types.all;
entity Comparator_1Bit_tb is
end Comparator_1Bit_tb;
