library verilog;
use verilog.vl_types.all;
entity Bh_FullAdder_tb is
end Bh_FullAdder_tb;
